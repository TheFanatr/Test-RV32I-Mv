`ifndef TYPES_SVH
`define TYPES_SVH
 
 

`endif // TYPES_SVH