`include "types.svh"

module rv32i (
    input clk,
    input clk_en,
    input rst
);

always @(posedge clk) begin
  //$display("CPU");
end

endmodule
