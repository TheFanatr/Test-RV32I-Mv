`timescale 1ns / 1ps

module core (
    input clk,
    input clk_en,
    input rst
);
    
endmodule